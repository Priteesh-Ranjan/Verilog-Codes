`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Institute: NIT Rourkela 
// Create Date: 13.01.2023 00:53:02
// Design Name: Priteesh Ranjan
// Module Name: Mux
// Project Name: 4x1 Mux 
//////////////////////////////////////////////////////////////////////////////////

module and_gate(a,b,c);
input a,b;
output c;
and(c,a,b);
endmodule
