`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Institute: NIT Rourkela 
// Create Date: 15.01.2023 00:20:39
// Design Name: Priteesh Ranjan
// Module Name: OR gate
// Project Name: orGate
//////////////////////////////////////////////////////////////////////////////////


module or_gate(a,b,c);
input a,b;
output c;
assign c = a|b;
endmodule
